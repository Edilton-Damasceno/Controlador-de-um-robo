module Robo (clock, reset, head, left, avancar, girar);


endmodule
